/*
    Jail Programming Language Copyright (C) 2022 SolindekDev

	Contribuitors:
		https://github.com/SolindekDev/Jail/edit/main/contributors.md
*/

module ast

// Enum of keywords
enum Keywords {
	puts = 0
	__rust
}

// String representation of enum
const (
	keyword_puts = "puts"
	keyword___rust = "__rust"
)
