module lexer

pub fn lexer() {
	println("Lexer")
}