module compiler

import os
import rand
import ast

pub fn str_to_byte(str string) []byte {
	mut bytes := []byte{}

	for i in str {
		bytes << i
	}	

	return bytes
}

fn writef(mut fs os.File, str string) {
	fs.write(
		str_to_byte(str)
	) or {
		println("cannot write to out.rs. not enough permissions.") 
		exit(1)
	}
}

pub fn compiler_init(mast ast.MainAST, out_flag bool) {
	mut out := os.create("out.rs") or {
		println("out.rs already exists")
		exit(1)
	}

	writef(mut out, "/*
    Jail Programming Language Copyright (C) 2022 SolindekDev
        - Code generated by Jail Programming Language
*/\n")
	writef(mut out, "
use std::io;
use std::process;\n")
	writef(mut out, "
#[warn(unused_variables)]
#[warn(unused_mut)]
#[warn(unused_imports)]
#[warn(unused_features)]
#[warn(dead_code)]
#[warn(non_snake_case)]
#[warn(non_upper_case_globals)]
#[warn(unreachable_code)]
#[warn(while_true)]
#[warn(unused_unsafe)]\n")
	writef(mut out, "
type int     = i32;
type uint    = i8;
type float   = f64;
type ufloat  = f32;\n")
	writef(mut out, "
fn main() {
")

	for i := 0; i < mast.body.len; i++ {
		actual_node_ast := mast.body[i]
		if actual_node_ast.type_ast == ast.TypeExpressionAST.ast_math_operation {
			body_tokens   := actual_node_ast.body_tokens
			mut operation := ""

			for j := 0; j < body_tokens.len; j++ {
				operation += body_tokens[j].value
			}

			name := rand.i64_in_range(0, 2000000)
			writef(mut out, "	let calculations_$name: float = ($operation) as float;\n")
		}		
	}
	writef(mut out, "}")

	out.close()

	os.execute("rustc out.rs")
	if out_flag == false { 
		os.execute("rm out.rs") 
	}
	os.execute("rm out.pdb")
}