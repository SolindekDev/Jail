module ast

enum Keywords {
	puts = 0
	exit
}

const (
	keyword_puts = "puts"
	keyword_exit = "exit"
)